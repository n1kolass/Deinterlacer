parameter DATA_WIDTH = 8;
parameter WIDTH = 640;
parameter HEIGHT = 480;
parameter HALF_HEIGHT = HEIGHT/2;